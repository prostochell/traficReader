module char_rom (
    input wire [7:0] char,    
    input wire [3:0] row,     
    output reg [7:0] data     
);


    reg [7:0] font [0:127][0:15];

    initial begin
		  // ASCII character '0' (0x30)
        font[8'h30][0]  = 8'b00111100;
        font[8'h30][1]  = 8'b01100110;
        font[8'h30][2]  = 8'b01101110;
        font[8'h30][3]  = 8'b01111110;
        font[8'h30][4]  = 8'b01110110;
        font[8'h30][5]  = 8'b01100110;
        font[8'h30][6]  = 8'b00111100;
        font[8'h30][7]  = 8'b00000000;
        font[8'h30][8]  = 8'b00000000;
        font[8'h30][9]  = 8'b00000000;
        font[8'h30][10] = 8'b00000000;
        font[8'h30][11] = 8'b00000000;
        font[8'h30][12] = 8'b00000000;
        font[8'h30][13] = 8'b00000000;
        font[8'h30][14] = 8'b00000000;
        font[8'h30][15] = 8'b00000000;

        // ASCII character '1' (0x31)
        font[8'h31][0]  = 8'b00011000;
        font[8'h31][1]  = 8'b00111000;
        font[8'h31][2]  = 8'b00011000;
        font[8'h31][3]  = 8'b00011000;
        font[8'h31][4]  = 8'b00011000;
        font[8'h31][5]  = 8'b00011000;
        font[8'h31][6]  = 8'b01111110;
        font[8'h31][7]  = 8'b00000000;
        font[8'h31][8]  = 8'b00000000;
        font[8'h31][9]  = 8'b00000000;
        font[8'h31][10] = 8'b00000000;
        font[8'h31][11] = 8'b00000000;
        font[8'h31][12] = 8'b00000000;
        font[8'h31][13] = 8'b00000000;
        font[8'h31][14] = 8'b00000000;
        font[8'h31][15] = 8'b00000000;

        // ASCII character '2' (0x32)
        font[8'h32][0]  = 8'b00111100;
        font[8'h32][1]  = 8'b01100110;
        font[8'h32][2]  = 8'b00000110;
        font[8'h32][3]  = 8'b00001100;
        font[8'h32][4]  = 8'b00110000;
        font[8'h32][5]  = 8'b01100000;
        font[8'h32][6]  = 8'b01111110;
        font[8'h32][7]  = 8'b00000000;
        font[8'h32][8]  = 8'b00000000;
        font[8'h32][9]  = 8'b00000000;
        font[8'h32][10] = 8'b00000000;
        font[8'h32][11] = 8'b00000000;
        font[8'h32][12] = 8'b00000000;
        font[8'h32][13] = 8'b00000000;
        font[8'h32][14] = 8'b00000000;
        font[8'h32][15] = 8'b00000000;

        // ASCII character '3' (0x33)
        font[8'h33][0]  = 8'b00111100;
        font[8'h33][1]  = 8'b01100110;
        font[8'h33][2]  = 8'b00000110;
        font[8'h33][3]  = 8'b00011100;
        font[8'h33][4]  = 8'b00000110;
        font[8'h33][5]  = 8'b01100110;
        font[8'h33][6]  = 8'b00111100;
        font[8'h33][7]  = 8'b00000000;
        font[8'h33][8]  = 8'b00000000;
        font[8'h33][9]  = 8'b00000000;
        font[8'h33][10] = 8'b00000000;
        font[8'h33][11] = 8'b00000000;
        font[8'h33][12] = 8'b00000000;
        font[8'h33][13] = 8'b00000000;
        font[8'h33][14] = 8'b00000000;
        font[8'h33][15] = 8'b00000000;

        // ASCII character '4' (0x34)
        font[8'h34][0]  = 8'b00001100;
        font[8'h34][1]  = 8'b00011100;
        font[8'h34][2]  = 8'b00111100;
        font[8'h34][3]  = 8'b01101100;
        font[8'h34][4]  = 8'b01111110;
        font[8'h34][5]  = 8'b00001100;
        font[8'h34][6]  = 8'b00001100;
        font[8'h34][7]  = 8'b00000000;
        font[8'h34][8]  = 8'b00000000;
        font[8'h34][9]  = 8'b00000000;
        font[8'h34][10] = 8'b00000000;
        font[8'h34][11] = 8'b00000000;
        font[8'h34][12] = 8'b00000000;
        font[8'h34][13] = 8'b00000000;
        font[8'h34][14] = 8'b00000000;
        font[8'h34][15] = 8'b00000000;

        // ASCII character '5' (0x35)
        font[8'h35][0]  = 8'b01111110;
        font[8'h35][1]  = 8'b01100000;
        font[8'h35][2]  = 8'b01111100;
        font[8'h35][3]  = 8'b00000110;
        font[8'h35][4]  = 8'b00000110;
        font[8'h35][5]  = 8'b01100110;
        font[8'h35][6]  = 8'b00111100;
        font[8'h35][7]  = 8'b00000000;
        font[8'h35][8]  = 8'b00000000;
        font[8'h35][9]  = 8'b00000000;
        font[8'h35][10] = 8'b00000000;
        font[8'h35][11] = 8'b00000000;
        font[8'h35][12] = 8'b00000000;
        font[8'h35][13] = 8'b00000000;
        font[8'h35][14] = 8'b00000000;
        font[8'h35][15] = 8'b00000000;

        // ASCII character '6' (0x36)
        font[8'h36][0]  = 8'b00111100;
        font[8'h36][1]  = 8'b01100110;
        font[8'h36][2]  = 8'b01100000;
        font[8'h36][3]  = 8'b01111100;
        font[8'h36][4]  = 8'b01100110;
        font[8'h36][5]  = 8'b01100110;
        font[8'h36][6]  = 8'b00111100;
        font[8'h36][7]  = 8'b00000000;
        font[8'h36][8]  = 8'b00000000;
        font[8'h36][9]  = 8'b00000000;
        font[8'h36][10] = 8'b00000000;
        font[8'h36][11] = 8'b00000000;
        font[8'h36][12] = 8'b00000000;
        font[8'h36][13] = 8'b00000000;
        font[8'h36][14] = 8'b00000000;
        font[8'h36][15] = 8'b00000000;

        // ASCII character '7' (0x37)
        font[8'h37][0]  = 8'b01111110;
        font[8'h37][1]  = 8'b00000110;
        font[8'h37][2]  = 8'b00001100;
        font[8'h37][3]  = 8'b00011000;
        font[8'h37][4]  = 8'b00110000;
        font[8'h37][5]  = 8'b01100000;
        font[8'h37][6]  = 8'b01100000;
        font[8'h37][7]  = 8'b00000000;
        font[8'h37][8]  = 8'b00000000;
        font[8'h37][9]  = 8'b00000000;
        font[8'h37][10] = 8'b00000000;
        font[8'h37][11] = 8'b00000000;
        font[8'h37][12] = 8'b00000000;
        font[8'h37][13] = 8'b00000000;
        font[8'h37][14] = 8'b00000000;
        font[8'h37][15] = 8'b00000000;

        // ASCII character '8' (0x38)
        font[8'h38][0]  = 8'b00111100;
        font[8'h38][1]  = 8'b01100110;
        font[8'h38][2]  = 8'b01100110;
        font[8'h38][3]  = 8'b00111100;
        font[8'h38][4]  = 8'b01100110;
        font[8'h38][5]  = 8'b01100110;
        font[8'h38][6]  = 8'b00111100;
        font[8'h38][7]  = 8'b00000000;
        font[8'h38][8]  = 8'b00000000;
        font[8'h38][9]  = 8'b00000000;
        font[8'h38][10] = 8'b00000000;
        font[8'h38][11] = 8'b00000000;
        font[8'h38][12] = 8'b00000000;
        font[8'h38][13] = 8'b00000000;
        font[8'h38][14] = 8'b00000000;
        font[8'h38][15] = 8'b00000000;

        // ASCII character '9' (0x39)
        font[8'h39][0]  = 8'b00111100;
        font[8'h39][1]  = 8'b01100110;
        font[8'h39][2]  = 8'b01100110;
        font[8'h39][3]  = 8'b00111110;
        font[8'h39][4]  = 8'b00000110;
        font[8'h39][5]  = 8'b01100110;
        font[8'h39][6]  = 8'b00111100;
        font[8'h39][7]  = 8'b00000000;
        font[8'h39][8]  = 8'b00000000;
        font[8'h39][9]  = 8'b00000000;
        font[8'h39][10] = 8'b00000000;
        font[8'h39][11] = 8'b00000000;
        font[8'h39][12] = 8'b00000000;
        font[8'h39][13] = 8'b00000000;
        font[8'h39][14] = 8'b00000000;
        font[8'h39][15] = 8'b00000000;

        // ASCII character 'A' (0x41)
        font[8'h41][0]  = 8'b00011000;
        font[8'h41][1]  = 8'b00100100;
        font[8'h41][2]  = 8'b01000010;
        font[8'h41][3]  = 8'b01000010;
        font[8'h41][4]  = 8'b01111110;
        font[8'h41][5]  = 8'b01000010;
        font[8'h41][6]  = 8'b01000010;
        font[8'h41][7]  = 8'b01000010;
        font[8'h41][8]  = 8'b00000000;
        font[8'h41][9]  = 8'b00000000;
        font[8'h41][10] = 8'b00000000;
        font[8'h41][11] = 8'b00000000;
        font[8'h41][12] = 8'b00000000;
        font[8'h41][13] = 8'b00000000;
        font[8'h41][14] = 8'b00000000;
        font[8'h41][15] = 8'b00000000;

        // ASCII character 'B' (0x42)
        font[8'h42][0]  = 8'b01111100;
        font[8'h42][1]  = 8'b01000010;
        font[8'h42][2]  = 8'b01000010;
        font[8'h42][3]  = 8'b01111100;
        font[8'h42][4]  = 8'b01000010;
        font[8'h42][5]  = 8'b01000010;
        font[8'h42][6]  = 8'b01111100;
        font[8'h42][7]  = 8'b00000000;
        font[8'h42][8]  = 8'b00000000;
        font[8'h42][9]  = 8'b00000000;
        font[8'h42][10] = 8'b00000000;
        font[8'h42][11] = 8'b00000000;
        font[8'h42][12] = 8'b00000000;
        font[8'h42][13] = 8'b00000000;
        font[8'h42][14] = 8'b00000000;
        font[8'h42][15] = 8'b00000000;

        // ASCII character 'C' (0x43)
        font[8'h43][0]  = 8'b00111100;
        font[8'h43][1]  = 8'b01100110;
        font[8'h43][2]  = 8'b01000000;
        font[8'h43][3]  = 8'b01000000;
        font[8'h43][4]  = 8'b01000000;
        font[8'h43][5]  = 8'b01100110;
        font[8'h43][6]  = 8'b00111100;
        font[8'h43][7]  = 8'b00000000;
        font[8'h43][8]  = 8'b00000000;
        font[8'h43][9]  = 8'b00000000;
        font[8'h43][10] = 8'b00000000;
        font[8'h43][11] = 8'b00000000;
        font[8'h43][12] = 8'b00000000;
        font[8'h43][13] = 8'b00000000;
        font[8'h43][14] = 8'b00000000;
        font[8'h43][15] = 8'b00000000;
		  
		  // ASCII character 'D' (0x44)
        font[8'h44][0]  = 8'b00000000;
        font[8'h44][1]  = 8'b00000000;
        font[8'h44][2]  = 8'b01111100;
        font[8'h44][3]  = 8'b01000010;
        font[8'h44][4]  = 8'b01000010;
        font[8'h44][5]  = 8'b01000010;
        font[8'h44][6]  = 8'b01000010;
        font[8'h44][7]  = 8'b01000010;
        font[8'h44][8]  = 8'b01000010;
        font[8'h44][9]  = 8'b01111100;
        font[8'h44][10] = 8'b00000000;
        font[8'h44][11] = 8'b00000000;
        font[8'h44][12] = 8'b00000000;
        font[8'h44][13] = 8'b00000000;
        font[8'h44][14] = 8'b00000000;
        font[8'h44][15] = 8'b00000000;

        // ASCII character 'E' (0x45)
        font[8'h45][0]  = 8'b00000000;
        font[8'h45][1]  = 8'b00000000;
        font[8'h45][2]  = 8'b01111110;
        font[8'h45][3]  = 8'b01000000;
        font[8'h45][4]  = 8'b01000000;
        font[8'h45][5]  = 8'b01111100;
        font[8'h45][6]  = 8'b01000000;
        font[8'h45][7]  = 8'b01000000;
        font[8'h45][8]  = 8'b01000000;
        font[8'h45][9]  = 8'b01111110;
        font[8'h45][10] = 8'b00000000;
        font[8'h45][11] = 8'b00000000;
        font[8'h45][12] = 8'b00000000;
        font[8'h45][13] = 8'b00000000;
        font[8'h45][14] = 8'b00000000;
        font[8'h45][15] = 8'b00000000;
		  
        // ASCII character 'F' (0x46)
        font[8'h45][0]  = 8'b00000000;
        font[8'h45][1]  = 8'b00000000;
        font[8'h45][2]  = 8'b01111110;
        font[8'h45][3]  = 8'b01000000;
        font[8'h45][4]  = 8'b01000000;
        font[8'h45][5]  = 8'b01111100;
        font[8'h45][6]  = 8'b01000000;
        font[8'h45][7]  = 8'b01000000;
        font[8'h45][8]  = 8'b01000000;
        font[8'h45][9]  = 8'b01000000;
        font[8'h45][10] = 8'b00000000;
        font[8'h45][11] = 8'b00000000;
        font[8'h45][12] = 8'b00000000;
        font[8'h45][13] = 8'b00000000;
        font[8'h45][14] = 8'b00000000;
        font[8'h45][15] = 8'b00000000;
    end

    always @(*) begin
        data = font[char][row];
    end
endmodule
